module PS2KeyboardMemory(
input logic clk,
input logic rst,

input logic [7:0]scanCode,
input logic scanCodeReady,

input logic [7:0]asciiKeyAddress,
output logic [31:0]asciiKeyValue
);

typedef enum logic [7:0] {
	sc_1_exclamation = 8'h16,
	sc_2_at = 8'h1E,
	sc_3_pound = 8'h26,
	sc_4_dollar = 8'h25,
	sc_5_percent = 8'h2E,
	sc_6_caret = 8'h36,
	sc_7_ampersand = 8'h3D,
	sc_8_asterisk = 8'h3E,
	sc_9_leftparenthesis = 8'h46,
	sc_0_rightparenthesis = 8'h45,
	sc_dash_underscore = 8'h4E,
	sc_plus_equals = 8'h55,
	sc_backspace = 8'h66,
	
	sc_tab = 8'h0D,
	sc_q_Q = 8'h15,
	sc_w_W = 8'h1D,
	sc_e_E = 8'h24,
	sc_r_R = 8'h2D,
	sc_t_T = 8'h2C,
	sc_y_Y = 8'h35,
	sc_u_U = 8'h3C,
	sc_i_I = 8'h43,
	sc_o_O = 8'h44,
	sc_p_P = 8'h4D,
	sc_leftbracket_leftcurly = 8'h54,
	sc_rightbracket_rightcurly = 8'h5B,
	sc_pipe_backslash = 8'h5D,
	
	sc_a_A = 8'h1C,
	sc_s_S = 8'h1B,
	sc_d_D = 8'h23,
	sc_f_F = 8'h2B,
	sc_g_G = 8'h34,
	sc_h_H = 8'h33,
	sc_j_J = 8'h3B,
	sc_k_K = 8'h42,
	sc_l_L = 8'h4B,
	sc_colon_semicolon = 8'h4C,
	sc_doublequote_singlequote = 8'h52,
	sc_enter = 8'h5A,
	
	sc_leftshift = 8'h12,
	sc_z_Z = 8'h1A,
	sc_x_X = 8'h22,
	sc_c_C = 8'h21,
	sc_v_V = 8'h2A,
	sc_b_B = 8'h32,
	sc_n_N = 8'h31,
	sc_m_M = 8'h3A,
	sc_lessthan_comma = 8'h41,
	sc_greaterthan_period = 8'h49,
	sc_questionmark_forwardslash = 8'h4A,
	sc_rightshift = 8'h59,
	
	sc_leftctrl = 8'h14,
	sc_leftalt = 8'h11,
	
	sc_space = 8'h29,
	
	// Extended
	// (Two bytes per key code)
	sce_rightalt = 8'h11,
	sce_rightctrl = 8'h14,
	
	sce_up = 8'h75,
	sce_down = 8'h72,
	sce_left = 8'h6B,
	sce_right = 8'h74
	
} ScanCodes;

typedef enum logic [7:0] {
	ascii_exclamation = 8'h21,
	ascii_doublequote = 8'h22,
	ascii_pound = 8'h23,
	ascii_dollarsign = 8'h24,
	ascii_percent = 8'h25,
	ascii_ampersand = 8'h26,
	ascii_singlequote = 8'h27,
	ascii_leftparenthesis = 8'h28,
	ascii_rightparenthesis = 8'h29,
	ascii_asterisk = 8'h2A,
	ascii_plus = 8'h2B,
	ascii_comma = 8'h2C,
	ascii_dash = 8'h2D,
	ascii_period = 8'h2E,
	ascii_forwardslash = 8'h2F,
	
	ascii_0 = 8'h30,
	ascii_1 = 8'h31,
	ascii_2 = 8'h32,
	ascii_3 = 8'h33,
	ascii_4 = 8'h34,
	ascii_5 = 8'h35,
	ascii_6 = 8'h36,
	ascii_7 = 8'h37,
	ascii_8 = 8'h38,
	ascii_9 = 8'h39,
	ascii_colon = 8'h3A,
	ascii_semicolon = 8'h3B,
	ascii_lessthan = 8'h3C,
	ascii_equals = 8'h3D,
	ascii_greaterthan = 8'h3E,
	ascii_questionmark = 8'h3F,
	ascii_at = 8'h40,
	ascii_A = 8'h41,
	ascii_B = 8'h42,
	ascii_C = 8'h43,
	ascii_D = 8'h44,
	ascii_E = 8'h45,
	ascii_F = 8'h46,
	ascii_G = 8'h47,
	ascii_H = 8'h48,
	ascii_I = 8'h49,
	ascii_J = 8'h4A,
	ascii_K = 8'h4B,
	ascii_L = 8'h4C,
	ascii_M = 8'h4D,
	ascii_N = 8'h4E,
	ascii_O = 8'h4F,
	ascii_P = 8'h50,
	ascii_Q = 8'h51,
	ascii_R = 8'h52,
	ascii_S = 8'h53,
	ascii_T = 8'h54,
	ascii_U = 8'h55,
	ascii_V = 8'h56,
	ascii_W = 8'h57,
	ascii_X = 8'h58,
	ascii_Y = 8'h59,
	ascii_Z = 8'h5A,
	ascii_leftbracket = 8'h5B,
	ascii_backslash = 8'h5C,
	ascii_rightbracket = 8'h5D,
	ascii_caret = 8'h5E,
	ascii_underscore = 8'h5F,
	
	ascii_backtick = 8'h60,
	ascii_a = 8'h61,
	ascii_b = 8'h62,
	ascii_c = 8'h63,
	ascii_d = 8'h64,
	ascii_e = 8'h65,
	ascii_f = 8'h66,
	ascii_g = 8'h67,
	ascii_h = 8'h68,
	ascii_i = 8'h69,
	ascii_j = 8'h6A,
	ascii_k = 8'h6B,
	ascii_l = 8'h6C,
	ascii_m = 8'h6D,
	ascii_n = 8'h6E,
	ascii_o = 8'h6F,
	ascii_p = 8'h70,
	ascii_q = 8'h71,
	ascii_r = 8'h72,
	ascii_s = 8'h73,
	ascii_t = 8'h74,
	ascii_u = 8'h75,
	ascii_v = 8'h76,
	ascii_w = 8'h77,
	ascii_x = 8'h78,
	ascii_y = 8'h79,
	ascii_z = 8'h7A,
	
	ascii_leftcurlybrace = 8'h7B,
	ascii_pipe = 8'h7C,
	ascii_rightcurlybrace = 8'h7D,
	ascii_tilde = 8'h7E,
	ascii_delete = 8'h7F
} AsciiCodes;


endmodule






