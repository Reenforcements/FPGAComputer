module RegisterFile_TB;


endmodule
