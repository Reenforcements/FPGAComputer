module LEDDisplayTest(
	input logic clk,
	input logic rst
);




endmodule