module PS2Keyboard_TB;

 logic clk;
 logic rst;

 logic PS2_CLK;
 logic PS2_DAT;

 logic [7:0]scanCode;
 logic scanCodeReady;
);


endmodule