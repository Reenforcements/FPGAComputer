module PS2KeyboardMemory_TB;




endmodule